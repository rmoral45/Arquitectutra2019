module rom
#(
    parameter NB_ROM_WORD   = 16,
    parameter NB_ROM_DEPTH  = 11,
    parameter DEPTH         = 2**NB_ROM_DEPTH
)
